//`ifndef b2gfifo_PKG_SV
//`define b2gfifo_PKG_SV

//------------------------------------------------------------------------------------------------------------
`include "uvm_macros.svh"

package b2gfifo_pkg;
    import uvm_pkg::*;
    
endpackage 

//`endif //b2gfifo_PKG_SV

