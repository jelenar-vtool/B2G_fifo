
//`include "uvm_pkg.sv"
`include "uvm_macros.svh" 
`include "b2gfifo_pkg.sv"
package b2gfifo_env_pkg;

import uvm_pkg::*;
import b2gfifo_pkg::*;


endpackage 

//------------------------------------------------------------------------------------------------------------


