class b2gfifo_cfg extends uvm_object;  

    // TODO: * * * Declare all the config fields * * *
    
    // TODO: * * * Register all the config fields with the factory* * *
    
    extern function new(string name = "b2gfifo_cfg");
    
    // TODO: * * * Define the set_default_config function * * *
endclass : b2gfifo_cfg

//-------------------------------------------------------------------------------------------------------------
function b2gfifo_cfg::new(string name = "b2gfifo_cfg");
    super.new(name);
endfunction : new


