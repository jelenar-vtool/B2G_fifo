`ifndef ENV_PKG_SV
`define ENV_PKG_SV

 `include "ahb_interface.sv"

package env_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "ahb_sequence_item.sv"
  `include "ahb_sequences.sv"
  `include "ahb_sequencer.sv"
  `include "ahb_driver.sv"
  `include "ahb_monitor.sv"
  `include "ahb_agent.sv"
  `include "ahb_scoreboard.sv"
  `include "ahb_environment.sv"

endpackage

`endif




