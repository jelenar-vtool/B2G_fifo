
//`include "uvm_pkg.sv"
`include "uvm_macros.svh" 
`include "temp_pkg.sv"
package temp_test_pkg;

import uvm_pkg::*;
import temp_pkg::*;

// * * * You can include different sequences for specific test bellow * * *

endpackage 

//------------------------------------------------------------------------------------------------------------


