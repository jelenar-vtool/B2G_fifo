`include "uvm_macros.svh" 
package fifo_ral_pkg;

import uvm_pkg::*;

endpackage 
