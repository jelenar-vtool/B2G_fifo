`include "uvm_macros.svh"
`include "env_pkg.sv"

module top;
    
    import uvm_pkg::*;
    import env_pkg::*;


endmodule
