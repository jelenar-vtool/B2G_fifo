`include "uvm_macros.svh"
`include "fifo_pkg.sv"
`include "fifo_ral_pkg.sv"

package fifo_env_pkg;

import uvm_pkg::*;
import fifo_pkg::*;
import fifo_ral_pkg::*;


endpackage 



