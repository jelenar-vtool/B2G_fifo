class b2gfifo_env_cfg extends uvm_object;       

    // TODO: * * * Declare all the env config fields * * *
    
    // TODO: * * * Declare all the lower-level config objects * * *

    // TODO: * * * Register all the config fields with the factory* * *

    extern function new(string name = "b2gfifo_env_cfg");
    
    // TODO: * * * Define the set_default_config function * * *
endclass

//-------------------------------------------------------------------------------------------------------------
function b2gfifo_env_cfg::new(string name = "b2gfifo_env_cfg");
    super.new(name);
    // TODO: * * * Instantiate the lower-level config objects * * *
endfunction
