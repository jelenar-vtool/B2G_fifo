
//`include "uvm_pkg.sv"
`include "uvm_macros.svh" 
`include "fifo_pkg.sv"
package fifo_test_pkg;

import uvm_pkg::*;
import fifo_pkg::*;

// * * * You can include different sequences for specific test bellow * * *

endpackage 

//------------------------------------------------------------------------------------------------------------


