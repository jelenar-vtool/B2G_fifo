`include "uvm_macros.svh" 
package ral_pkg;

import uvm_pkg::*;

endpackage 
