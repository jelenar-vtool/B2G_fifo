
`include "b2gfifo_base_test.sv"
`include "b2gfifo_extended_test.sv"
`include "b2gfifo_random_test.sv"            
`include "b2gfifo_rst_test.sv"
