
//`include "uvm_pkg.sv"

package b2gfifo_test_pkg;

    import uvm_pkg::*;
    import b2gfifo_pkg::*;
    import b2gfifo_env_pkg::*;
    
    `include "uvm_macros.svh" 
    `include "b2gfifo_base_test.sv"

    // * * * You can include different sequences for specific test bellow * * *

endpackage 

//------------------------------------------------------------------------------------------------------------


