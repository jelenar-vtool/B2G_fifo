`timescale 1ns/100ps

parameter bit [5:0] go_duration = 50;
parameter bit [5:0] go_stop_duration = 5;
parameter bit [5:0] stop_duration = 20;
parameter bit [5:0] stop_go_duration = 2;

parameter daytime   = 1'b0;
parameter nighttime = 1'b1;
parameter go = 2'b00;
parameter go_stop = 2'b01;
parameter stop = 2'b10;
parameter stop_go = 2'b11;

module traffic_lights (
	input logic clk,
	input logic rst_n,
	input logic broken,
	output logic r_l,
	output logic y_l,
	output logic g_l
);
	
	parameter bit [9:0] day_duration = 600;
	parameter bit [9:0] night_duration = 200;

	enum bit {DAYTIME, NIGHTTIME} time_of_day;
	enum bit [1:0] {GO, GO_STOP, STOP, STOP_GO} lights_state;

	bit yellow_on;

	bit Q, nextQ;
	bit [1:0] QQ, nextQQ;
	bit day_switch;
	bit lights_switch;

	bit [9:0] day_switch_cnt = 0;
	bit [9:0] day_switch_cnt_th = day_duration;

	bit [5:0] lights_switch_cnt = 0;
	bit [5:0] lights_switch_cnt_th = go_duration;


	// ----------------------------------------------------------------------
	// EXERCISE 4
	// a) Comment out line with `include statement, which is BELOW
	//    and run the simulation. It will reveal the bug in RTL.
	// b) Find this bug based on the errors generated by blinking 
	//    yellow light assertion from exercise 3
	// If you find it, it means you are a real PRO in a BUG HUNTING WORLD :D
	// ----------------------------------------------------------------------
	// YOUR CODE HERE - START
	








	// YOUR CODE HERE - END
	// ----------------------------------------------------------------------
	`include "solutions/ex4_solved.v"

	// Current state register
	always @(posedge clk) begin
		if(rst_n) begin
			nextQ = DAYTIME;
			nextQQ = GO;
		end
		else begin
			Q = nextQ;
			QQ = nextQQ;
		end
	end

	// Day - Night counter
	always @(posedge clk) begin
		if(rst_n) begin
			day_switch_cnt = 0;
			day_switch = 0;
		end

		day_switch_cnt = day_switch_cnt + 1'b1;
		day_switch = 0;

		if (day_switch_cnt == day_switch_cnt_th) begin
			day_switch_cnt = 0;
			day_switch = 1;
		end
	end

	// Lights counter
	always @(posedge clk) begin
		if(rst_n) begin
			lights_switch_cnt = 0;
			lights_switch = 0;
		end

		lights_switch_cnt = lights_switch_cnt + 1'b1;
		lights_switch = 0;

		if (lights_switch_cnt == lights_switch_cnt_th) begin
			lights_switch_cnt = 0;
			lights_switch = 1;
		end
	end


	// Day - Night logic
	always @(posedge clk) begin
		nextQ = 1'bx;
		case(Q)
		DAYTIME:
			if(day_switch) begin
				time_of_day = NIGHTTIME; 
				day_switch_cnt_th = night_duration;
			end
			else begin			
				time_of_day = DAYTIME;
			end
		NIGHTTIME:
			if(day_switch)	begin			
				time_of_day = DAYTIME;
				day_switch_cnt_th = day_duration;
			end
			else begin
				time_of_day = NIGHTTIME; 
			end
		endcase
		nextQ = time_of_day;
	end

	// Lights state logic
	always @(QQ or lights_switch) begin
		nextQQ = 2'bxx;
		case(QQ)
		GO:
			if(lights_switch) begin
				lights_state = GO_STOP;
				lights_switch_cnt_th = go_stop_duration;
			end
			else begin
				lights_state = GO;
			end
		GO_STOP:
			if(lights_switch) begin
				lights_state = STOP;
				lights_switch_cnt_th = stop_duration;
			end
			else begin
				lights_state = GO_STOP;
			end
		STOP:
			if(lights_switch) begin
				lights_state = STOP_GO;
				lights_switch_cnt_th = stop_go_duration;
			end
			else begin
				lights_state = STOP;
			end
		STOP_GO:
			if(lights_switch) begin
				lights_state = GO;
				lights_switch_cnt_th = go_duration;
			end
			else begin
				lights_state = STOP_GO;
			end
		endcase
		nextQQ = lights_state;
	end

	always @(posedge clk) begin
		if (nextQ == NIGHTTIME)
			yellow_on = ~yellow_on;
	end

	// always @(posedge clk or Q or QQ) begin
	always @(posedge clk) begin
		r_l = 0;
		y_l = 0;
		g_l = 0;

		case(Q)
		DAYTIME: begin
			case(QQ)
			GO: begin
				r_l = 0;
				y_l = 0;
				g_l = 1;
			end
			GO_STOP: begin
				r_l = 0;
				y_l = 1;
				g_l = 0;
			end
			STOP: begin
				r_l = 1;
				y_l = 0;
				g_l = 0;
			end	
			STOP_GO: begin
				r_l = 1;
				y_l = 1;
				g_l = 0;
			end
			endcase
		end
		NIGHTTIME:
			if(yellow_on) begin
				r_l = 0;
				y_l = 1;
				g_l = 0;
			end
			else begin //YELLOW_OFF
				r_l = 0;
				y_l = 0;
				g_l = 0;
			end
		endcase
	end

	task wait_clk (input int no_clocks);
	begin
		repeat (no_clocks) @ (posedge clk);
	end
	endtask


endmodule //DUT
