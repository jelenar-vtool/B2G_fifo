class b2gfifo_virtual_sequencer extends uvm_sequencer #(b2gfifo_item);
    // TODO: * * * Declare the sequencer handle * * *
    
    // TODO: * * * Add to factory * * *

    // TODO: * * * Declare and define other necessary tasks and functions * * *
endclass : b2gfifo_virtual_sequencer
