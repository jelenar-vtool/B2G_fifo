
//`include "uvm_pkg.sv"
`include "uvm_macros.svh" 
`include "b2gfifo_pkg.sv"
package b2gfifo_test_pkg;

import uvm_pkg::*;
    import b2gfifo_pkg::*;

    `include "b2gfifo_simple_base_test.sv"

// * * * You can include different sequences for specific test bellow * * *

endpackage 

//------------------------------------------------------------------------------------------------------------


