`include "uvm_macros.svh"
`include "fifo_env_pkg.sv"

module top;
    
    import uvm_pkg::*;
    import fifo_env_pkg::*;


endmodule
