`include "uvm_macros.svh"
`include "uvc_pkg.sv"

package env_pkg;

import uvm_pkg::*;
import uvc_pkg::*;


endpackage 



