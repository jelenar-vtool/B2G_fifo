//------------------------------------------------------------------------------------------------------------
package b2gfifo_env_pkg;
    import uvm_pkg::*;
    import b2gfifo_pkg::*;

   //`include "b2gfifo_cfg.sv"
   `include "b2gfifo_virtual_sequencer.sv"
   //`include "b2gfifo_agent.sv" 
   `include "b2gfifo_env_cfg.sv"
   `include "b2gfifo_scoreboard.sv"

   `include "b2gfifo_virtual_sequence.sv"
   `include "b2gfifo_env.sv"

endpackage 

//------------------------------------------------------------------------------------------------------------


