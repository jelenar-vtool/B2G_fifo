`include "uvm_macros.svh" 

package b2gfifo_test_pkg;

    import uvm_pkg::*;
    import b2gfifo_pkg::*;
    import b2gfifo_env_pkg::*;

    `include "b2gfifo_simple_base_test.sv"
endpackage 
