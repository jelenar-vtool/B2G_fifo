
interface b2gfifo_if;
    // * * * TODO: Add all the necessary interface signals and logic * * *

endinterface   
    


