
interface b2gfifo_topvif();
  logic clk;
  logic rst_n;

  //Declare all inputs and outputs



endinterface
  
