//------------------------------------------------------------------------------------------------------------
package b2gfifo_env_pkg;
    import uvm_pkg::*;
    import b2gfifo_pkg::*;
    
    `include "uvm_macros.svh" 
    `include "b2gfifo_env_cfg.sv"
    `include "b2gfifo_env.sv"
endpackage 
