
`include "fifo_base_test.sv"
