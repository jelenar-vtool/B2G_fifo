`ifndef TEST_PKG_SV
`define TEST_PKG_SV


package test_lib_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import env_pkg::*;

  `include "ahb_base_test.sv"
  `include "ahb_write_read_test.sv"

endpackage

`endif


