// TODO: * * * Write the extended test class here * * *

// TODO: * * * Extend this class from base test class * * *

// TODO: * * * Add to factory and declare a virtual sequence for this test * * *

// TODO: * * * Declare the test constructor and run_phase task * * *

// TODO: * * * Write the test constructor definition * * *

// TODO: * * * Write the run_phase definition. Randomize and start the virtual sequence in it * * *

// TODO: * * * Don't forget to add the objections! * * *
