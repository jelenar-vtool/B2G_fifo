
`include "temp_base_test.sv"
`include "temp_extended_test.sv"
`include "temp_random_test.sv"            
`include "temp_rst_test.sv"
