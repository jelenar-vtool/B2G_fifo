
interface fifo_if (input bit system_clock, input bit reset_n);
    
    // * * * Add you specific interface logics below * * *

    // * * * You can add assertion checkers bellow * * * 
    

endinterface   
    


