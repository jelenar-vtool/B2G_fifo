`include "uvm_macros.svh"

package uvc_pkg;

import uvm_pkg::*;


endpackage 



