`include "uvm_macros.svh"

package fifo_pkg;

import uvm_pkg::*;


endpackage 



